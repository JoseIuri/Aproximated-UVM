`ifndef MUL8S_TYPES
`define MUL8S_TYPES

`endif